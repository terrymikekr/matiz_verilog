module m2(
input d,
input e,

output f


);



m1 m3(
.a(d),
.b(e),
.c(f)
);



endmodule
